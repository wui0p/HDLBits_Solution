module top_module(output zero);
    //this module does not need any code
    //wire is automatically set to 0 in Verilog
endmodule
