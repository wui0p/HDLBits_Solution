module top_module (
    output out);

    //all variable is set to 0 as default
    //thus a GND wire do not have to do anything

endmodule