module top_module (
    input in,
    output out);

    //connect 'in' wire to 'out', using assign
    assign out = in;
    
endmodule