module top_module( input in, output out );

    //connecting wire output to wire input 
    assign out = in;
    
endmodule