module top_module( output one );

    //this assign wire "one" as 1, infinitly
    assign one = 1;

endmodule