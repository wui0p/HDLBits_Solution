module top_module( input in, output out );

    // '~' or '!' work as NOT gate
    assign out = ~in;
    
endmodule